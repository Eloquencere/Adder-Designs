class adder_test_config extends uvm_object;
    `uvm_object_utils(adder_test_config)

    function new(string name = "adder_test_config");
        super.new(name);
    endfunction
endclass
