class packet;
    randc bit [15:0]a, b;
    randc bit cin;
    bit [15:0]sum;
    bit cout;
endclass
