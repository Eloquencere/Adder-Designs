module pipline (

);

endmodule
