`timescale 1ns / 1ps

interface DUT_interface();
    logic [15:0]a,b;
    logic cin;
    logic [15:0]sum;
    logic cout;
endinterface
