package adder_sequences_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "sequence_item/adder_sequence_item.sv"
	
	`include "basic_operation_sequence.sv"
	`include "single_bit_sequence.sv"
	`include "zero_propagation_sequence.sv"
	`include "carry_propagation_sequence.sv"
	`include "overflow_sequence.sv"
	`include "underflow_sequence.sv"
	`include "random_no_constraint_sequence.sv"
endpackage