package adder_testbench_constants_pkg;
    parameter bit colourise_report_message = 1;

    parameter string dut_list[] = '{
        "CIAxbit"
        // "CLAxbit",
        // "CSelAxbit",
        // "CSkAxbit",
        // "RCAxbit",
        // "MCCAxbit"
    };
endpackage


