package adder_testbench_constants_pkg;
    parameter string dut_list[] = 
    {
        "CIAxbit",
        "CLAxbit",
        "CSelAxbit",
        "CSkAxbit",
        "RCAxbit",
        "MCCAxbit"
    };
endpackage
